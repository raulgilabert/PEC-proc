LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE IEEE.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY Tarea8 IS
	PORT( CLOCK_50 : IN std_logic;
			HEX0 : OUT std_logic_vector(6 downto 0);
			HEX1 : OUT std_logic_vector(6 downto 0);
			HEX2 : OUT std_logic_vector(6 downto 0);
			HEX3 : OUT std_logic_vector(6 downto 0));
END Tarea8;

ARCHITECTURE Structure OF Tarea8 IS
BEGIN
.
. -- Aquí debéis poner vuestro código que implemente la tarea
.
END Structure;